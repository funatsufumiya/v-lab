module main

import sub

fn main(){
	println("hello")
	sub.sub()
}