module main

fn main(){
	println("hello from V!")
}